module ucode_rom(
    output reg [34:0] control_store [0:63]
);
    initial begin
        control_store[0]  = 35'b01001001000000000000000000000000000;
        control_store[1]  = 35'b00001001000001100010000010000000000;
        control_store[2]  = 35'b00001110110000000001000011011000000;
        control_store[3]  = 35'b00001100010000000001000011011000000;
        control_store[4]  = 35'b01101010000000000000000000000000000;
        control_store[5]  = 35'b00001001000001100010000010000010000;
        control_store[6]  = 35'b00001100110000000001000011011000001;
        control_store[7]  = 35'b00001011110000000001000011011000001;
        control_store[8]  = 35'b00000000000000000000000000000000000;
        control_store[9]  = 35'b00001001000001100010000010000100000;
        control_store[10] = 35'b00000000000000000000000000000000000;
        control_store[11] = 35'b00000000000000000000000000000000000;
        control_store[12] = 35'b00001001000000010000010011000000000;
        control_store[13] = 35'b00001001000001100000100010000000000;
        control_store[14] = 35'b00001001000001000001000000101000001;
        control_store[15] = 35'b00001110010000000001000000000000000;
        control_store[16] = 35'b00101000000000000000000000000001110;
        control_store[17] = 35'b00101000100000000000000000000001100;
        control_store[18] = 35'b00010000110000011000000000001000000;
        control_store[19] = 35'b00010000110000011000000000001000000;
        control_store[20] = 35'b00001001000001011000010111000000000;
        control_store[21] = 35'b00001001000001011000010100110000001;
        control_store[22] = 35'b00001001000000010000010000100000001;
        control_store[23] = 35'b00001000001000000010000000000110010;
        control_store[24] = 35'b00001000101000000010000000000110000;
        control_store[25] = 35'b00101100101000000000000000000001010;
        control_store[26] = 35'b00000000000000000000000000000000000;
        control_store[27] = 35'b00001001000001100100000000000000010;
        control_store[28] = 35'b00101110001001001000000100000001010;
        control_store[29] = 35'b00101110101000000000000000000001000;
        control_store[30] = 35'b00001001000000010100001000000000010;
        control_store[31] = 35'b00001001000001100100000000000000000;
        control_store[32] = 35'b10000000000010000000000000000000000;
        control_store[33] = 35'b00110000101000000000000000000001010;
        control_store[34] = 35'b00000000000000000000000000000000000;
        control_store[35] = 35'b00010000000100000100000000000000010;
        control_store[36] = 35'b00000000000000000000000000000000000;
        control_store[37] = 35'b00000000000000000000000000000000000;
        control_store[38] = 35'b00000000000000000000000000000000000;
        control_store[39] = 35'b00000000000000000000000000000000000;
        control_store[40] = 35'b00000000000000000000000000000000000;
        control_store[41] = 35'b00000000000000000000000000000000000;
        control_store[42] = 35'b00000000000000000000000000000000000;
        control_store[43] = 35'b00000000000000000000000000000000000;
        control_store[44] = 35'b00000000000000000000000000000000000;
        control_store[45] = 35'b00000000000000000000000000000000000;
        control_store[46] = 35'b00000000000000000000000000000000000;
        control_store[47] = 35'b00000000000000000000000000000000000;
        control_store[48] = 35'b00000000000000000000000000000000000;
        control_store[49] = 35'b00000000000000000000000000000000000;
        control_store[50] = 35'b00000000000000000000000000000000000;
        control_store[51] = 35'b00000000000000000000000000000000000;
        control_store[52] = 35'b00000000000000000000000000000000000;
        control_store[53] = 35'b00000000000000000000000000000000000;
        control_store[54] = 35'b00000000000000000000000000000000000;
        control_store[55] = 35'b00000000000000000000000000000000000;
        control_store[56] = 35'b00000000000000000000000000000000000;
        control_store[57] = 35'b00000000000000000000000000000000000;
        control_store[58] = 35'b00000000000000000000000000000000000;
        control_store[59] = 35'b00000000000000000000000000000000000;
        control_store[60] = 35'b00000000000000000000000000000000000;
        control_store[61] = 35'b00000000000000000000000000000000000;
        control_store[62] = 35'b00000000000000000000000000000000000;
        control_store[63] = 35'b00000000000000000000000000000000000;
    end
endmodule