module ucode_rom();
endmodule