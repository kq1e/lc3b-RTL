module microsequencer();

endmodule