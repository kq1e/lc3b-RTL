module memory();
    input [15:0] ADDR,
    input 

endmodule