module LC3B_top(
    input CLK
);
    
    reg [15:0] PC;
    reg [15:0] IR;
endmodule
