module microsequencer();

endmodule

